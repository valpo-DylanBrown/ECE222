library ieee;
use ieee.std_logic_1164.all;

entity Elevator is
  port( );
end Elevator;

architecture behav of Elevator is

  signal

begin

end behav;
