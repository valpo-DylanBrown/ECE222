library ieee;
use ieee.std_logic_1164.all;

entity Elevator is
  port( );
end Elevator;

architecture behav of Elevator is
  type State is (S0, S1, S2, S3);
  signal

begin

end behav;
